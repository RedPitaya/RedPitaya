package str_pkg;

typedef struct {
  real fix;
  real rnd;
} tmg_t;

endpackage: str_pkg
