////////////////////////////////////////////////////////////////////////////////
// Module: RLE (Run Length Encoding) compression
// Author: Iztok Jeras
// (c) Red Pitaya  http://www.redpitaya.com
////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////
//
// GENERAL DESCRIPTION:
//
// A RLE compression is applied to the signal.
////////////////////////////////////////////////////////////////////////////////

module rle #(
  // counter properties
  int unsigned CW = 8,
  // stream properties
  int unsigned DN = 1,
  type DTI = logic [8-1:0], // data type for input
  type DTO = logic [8-1:0]  // data type for output
)(
  // input stream input/output
  axi4_stream_if.d sti,  // input
  axi4_stream_if.s sto,  // output
  // configuration
  input  logic     ctl_rst,  // reset
  input  logic     cfg_ena   // enable
);

////////////////////////////////////////////////////////////////////////////////
// store previous value
////////////////////////////////////////////////////////////////////////////////

DTI   old_tdata ;
logic old_tvalid;
logic old_tlast ;

always_ff @(posedge sti.ACLK)
if (sti.transf) begin
  old_tdata <= sti.TDATA;
  old_tlast <= sti.TLAST;
end

always_ff @(posedge sti.ACLK)
if (~sti.ARESETn)     old_tvalid <= 1'b0;
else if (sti.transf)  old_tvalid <= ~sti.TLAST;

////////////////////////////////////////////////////////////////////////////////
// comparator
////////////////////////////////////////////////////////////////////////////////

logic cmp;  // compare

assign cmp = (old_tdata == sti.TDATA);

////////////////////////////////////////////////////////////////////////////////
// counter
////////////////////////////////////////////////////////////////////////////////

logic [CW-1:0] cnt;
logic [CW-1:0] nxt;

always_ff @(posedge sti.ACLK)
if (~sti.ARESETn)     cnt <= '0;
else if (sti.transf)  cnt <= nxt;

assign nxt = cnt + 1;

////////////////////////////////////////////////////////////////////////////////
// output
////////////////////////////////////////////////////////////////////////////////

always_ff @(posedge sti.ACLK)
if (sti.transf)  sto.TLAST <= old_tlast;

assign sto.TDATA = {cnt, old_tdata};

endmodule: rle
