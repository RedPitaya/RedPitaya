////////////////////////////////////////////////////////////////////////////////
// Module: Red Pitaya TOP package.
// Authors: Iztok Jeras
// (c) Red Pitaya  http://www.redpitaya.com
////////////////////////////////////////////////////////////////////////////////

package top_pkg;

// module numbers
localparam int unsigned MNO = 2;  // number of oscilloscope modules
localparam int unsigned MNG = 2;  // number of generator    modules

// all events
typedef struct packed {
  osc_pkg::evn_t           la;   // logic analyzer
  gen_pkg::evn_t           lg;   // logic generator
  osc_pkg::evn_t [MNO-1:0] osc;  // oscilloscope
  gen_pkg::evn_t [MNG-1:0] gen;  // generator
} evn_t;

// interrupts
typedef struct packed {
  logic           la;   // logic analyzer
  logic           lg;   // logic generator
  logic [MNO-1:0] osc;  // oscilloscope
  logic [MNG-1:0] gen;  // generator
} irq_t;

endpackage: top_pkg
