////////////////////////////////////////////////////////////////////////////////
// Module: RLE (Run Length Encoding) compression
// Author: Iztok Jeras
// (c) Red Pitaya  http://www.redpitaya.com
////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////
//
// GENERAL DESCRIPTION:
//
// A RLE compression is applied to the signal.
//
////////////////////////////////////////////////////////////////////////////////

module rle #(
  // counter properties
  int unsigned CW = 8,
  // stream properties
  int unsigned DN = 1,
  type DTI = logic [8-1:0], // data type for input
  type DTO = logic [8-1:0]  // data type for output
)(
  // input stream input/output
  axi4_stream_if.d sti,  // input
  axi4_stream_if.s sto,  // output
  // configuration
  input  logic     ctl_rst,  // reset
  input  logic     cfg_ena   // enable
);

////////////////////////////////////////////////////////////////////////////////
// local variables
////////////////////////////////////////////////////////////////////////////////

// old values
DTI   old_tdata ;
logic old_tvalid;

// comparator
logic cmp;

// counter
logic [CW-1:0] cnt;
logic [CW-1:0] nxt;
logic          max;

// compression
logic trn;

////////////////////////////////////////////////////////////////////////////////
// store previous value
////////////////////////////////////////////////////////////////////////////////

always_ff @(posedge sti.ACLK)
if (sti.transf) begin
  old_tdata <= sti.TDATA;
end

always_ff @(posedge sti.ACLK)
if (~sti.ARESETn)     old_tvalid <= 1'b0;
else if (sti.transf)  old_tvalid <= ~sti.TLAST;

////////////////////////////////////////////////////////////////////////////////
// comparator
////////////////////////////////////////////////////////////////////////////////

assign cmp = (old_tdata == sti.TDATA);

////////////////////////////////////////////////////////////////////////////////
// counter
////////////////////////////////////////////////////////////////////////////////

assign nxt = cnt + 1;
assign max = &cnt;

always_ff @(posedge sti.ACLK)
if (~sti.ARESETn)     cnt <= '0;
else if (sti.transf)  cnt <= trn ? '0 : nxt;

////////////////////////////////////////////////////////////////////////////////
// compression
////////////////////////////////////////////////////////////////////////////////

assign trn = ~old_tvalid | ~cmp | max | sti.TLAST; 

assign sti.TREADY = sto.TREADY | ~sto.TVALID;

always_ff @(posedge sti.ACLK)
if (~sti.ARESETn)     sto.TVALID <= 1'b0;
else if (sti.transf)  sto.TVALID <= trn;

always_ff @(posedge sti.ACLK)
if (sti.transf) begin
  sto.TLAST <= sti.TLAST;
  sto.TKEEP <= sti.TKEEP;
end

assign sto.TDATA = {cnt, old_tdata};

endmodule: rle
