////////////////////////////////////////////////////////////////////////////////
// @brief Red Pitaya Processing System (PS) wrapper. Including simple AXI slave.
// @Author Matej Oblak
// (c) Red Pitaya  http://www.redpitaya.com
////////////////////////////////////////////////////////////////////////////////

/**
 * GENERAL DESCRIPTION:
 *
 * Wrapper of block design.  
 *
 *                   /-------\
 *   PS CLK -------> |       | <---------------------> SPI master & slave
 *   PS RST -------> |  PS   |
 *                   |       | ------------+---------> FCLK & reset 
 *                   |       |             |
 *   PS DDR <------> |  ARM  |   AXI   /-------\
 *   PS MIO <------> |       | <-----> |  AXI  | <---> system bus
 *                   \-------/         | SLAVE |
 *                                     \-------/
 *
 * Module wrappes PS module (BD design from Vivado or EDK from PlanAhead).
 * There is also included simple AXI slave which serves as master for custom
 * system bus. With this simpler bus it is more easy for newbies to develop 
 * their own module communication with ARM.
 */

module red_pitaya_ps (
  // PS peripherals
  inout  logic [ 54-1:0] FIXED_IO_mio       ,
  inout  logic           FIXED_IO_ps_clk    ,
  inout  logic           FIXED_IO_ps_porb   ,
  inout  logic           FIXED_IO_ps_srstb  ,
  inout  logic           FIXED_IO_ddr_vrn   ,
  inout  logic           FIXED_IO_ddr_vrp   ,
  // DDR
  inout  logic [ 15-1:0] DDR_addr           ,
  inout  logic [  3-1:0] DDR_ba             ,
  inout  logic           DDR_cas_n          ,
  inout  logic           DDR_ck_n           ,
  inout  logic           DDR_ck_p           ,
  inout  logic           DDR_cke            ,
  inout  logic           DDR_cs_n           ,
  inout  logic [  4-1:0] DDR_dm             ,
  inout  logic [ 32-1:0] DDR_dq             ,
  inout  logic [  4-1:0] DDR_dqs_n          ,
  inout  logic [  4-1:0] DDR_dqs_p          ,
  inout  logic           DDR_odt            ,
  inout  logic           DDR_ras_n          ,
  inout  logic           DDR_reset_n        ,
  inout  logic           DDR_we_n           ,
  // system signals
  input  logic           clk                ,
  input  logic           rstn               ,
  output logic [  4-1:0] fclk_clk_o         ,
  output logic [  4-1:0] fclk_rstn_o        ,
  // XADC
  input  logic  [ 5-1:0] vinp_i             ,  // voltages p
  input  logic  [ 5-1:0] vinn_i             ,  // voltages n
  // system read/write channel
  sys_bus_if.m           bus,
  axi4_lite_if.m         axi4_lite,
  // stream input
  str_bus_if.d           sti [2-1:0]
);

////////////////////////////////////////////////////////////////////////////////
// AXI SLAVE
////////////////////////////////////////////////////////////////////////////////

logic [4-1:0] fclk_clk ;
logic [4-1:0] fclk_rstn;

axi_bus_if #(.DW (32), .AW (32), .IW (12), .LW (4)) axi_gp (.ACLK (bus.clk), .ARESETn (rstn));

/*
axi_slave #(
  .DW (32),
  .AW (32),
  .IW (12)
) axi_slave_gp0 (
  // AXI bus
  .axi       (axi_gp),
  // system read/write channel
  .bus       (bus)
);
*/

axi4_slave_old #(
  .AXI_DW     (  32     ), // data width (8,16,...,1024)
  .AXI_AW     (  32     ), // address width
  .AXI_IW     (  12     )  // ID width
) axi_slave_gp0 (
  // global signals
  .axi_clk_i        (  axi_gp.ACLK           ),  // global clock
  .axi_rstn_i       (  rstn                  ),  // global reset
  // axi write address channel
  .axi_awid_i       (  axi_gp.AWID           ),  // write address ID
  .axi_awaddr_i     (  axi_gp.AWADDR         ),  // write address
  .axi_awlen_i      (  axi_gp.AWLEN          ),  // write burst length
  .axi_awsize_i     (  axi_gp.AWSIZE         ),  // write burst size
  .axi_awburst_i    (  axi_gp.AWBURST        ),  // write burst type
  .axi_awlock_i     (  axi_gp.AWLOCK         ),  // write lock type
  .axi_awcache_i    (  axi_gp.AWCACHE        ),  // write cache type
  .axi_awprot_i     (  axi_gp.AWPROT         ),  // write protection type
  .axi_awvalid_i    (  axi_gp.AWVALID        ),  // write address valid
  .axi_awready_o    (  axi_gp.AWREADY        ),  // write ready
  // axi write data channel
  .axi_wid_i        (  axi_gp.WID            ),  // write data ID
  .axi_wdata_i      (  axi_gp.WDATA          ),  // write data
  .axi_wstrb_i      (  axi_gp.WSTRB          ),  // write strobes
  .axi_wlast_i      (  axi_gp.WLAST          ),  // write last
  .axi_wvalid_i     (  axi_gp.WVALID         ),  // write valid
  .axi_wready_o     (  axi_gp.WREADY         ),  // write ready
  // axi write response channeL
  .axi_bid_o        (  axi_gp.BID            ),  // write response ID
  .axi_bresp_o      (  axi_gp.BRESP          ),  // write response
  .axi_bvalid_o     (  axi_gp.BVALID         ),  // write response valid
  .axi_bready_i     (  axi_gp.BREADY         ),  // write response ready
  // axi read address channel
  .axi_arid_i       (  axi_gp.ARID           ),  // read address ID
  .axi_araddr_i     (  axi_gp.ARADDR         ),  // read address
  .axi_arlen_i      (  axi_gp.ARLEN          ),  // read burst length
  .axi_arsize_i     (  axi_gp.ARSIZE         ),  // read burst size
  .axi_arburst_i    (  axi_gp.ARBURST        ),  // read burst type
  .axi_arlock_i     (  axi_gp.ARLOCK         ),  // read lock type
  .axi_arcache_i    (  axi_gp.ARCACHE        ),  // read cache type
  .axi_arprot_i     (  axi_gp.ARPROT         ),  // read protection type
  .axi_arvalid_i    (  axi_gp.ARVALID        ),  // read address valid
  .axi_arready_o    (  axi_gp.ARREADY        ),  // read address ready
  // axi read data channel
  .axi_rid_o        (  axi_gp.RID            ),  // read response ID
  .axi_rdata_o      (  axi_gp.RDATA          ),  // read data
  .axi_rresp_o      (  axi_gp.RRESP          ),  // read response
  .axi_rlast_o      (  axi_gp.RLAST          ),  // read last
  .axi_rvalid_o     (  axi_gp.RVALID         ),  // read response valid
  .axi_rready_i     (  axi_gp.RREADY         ),  // read response ready
  // system read/write channel
  .sys_addr_o       (  bus.addr              ),  // system read/write address
  .sys_wdata_o      (  bus.wdata             ),  // system write data
  .sys_sel_o        (                        ),  // system write byte select
  .sys_wen_o        (  bus.wen               ),  // system write enable
  .sys_ren_o        (  bus.ren               ),  // system read enable
  .sys_rdata_i      (  bus.rdata             ),  // system read data
  .sys_err_i        (  bus.err               ),  // system error indicator
  .sys_ack_i        (  bus.ack               )   // system acknowledge signal
);

//always @(posedge bus.clk)
//rstn <= fclk_rstn[0];

////////////////////////////////////////////////////////////////////////////////
// PS STUB
////////////////////////////////////////////////////////////////////////////////

assign fclk_rstn_o = fclk_rstn;

BUFG fclk_buf [4-1:0] (.O(fclk_clk_o), .I(fclk_clk));

system_wrapper system_i (
  // MIO
  .FIXED_IO_mio      (FIXED_IO_mio     ),
  .FIXED_IO_ps_clk   (FIXED_IO_ps_clk  ),
  .FIXED_IO_ps_porb  (FIXED_IO_ps_porb ),
  .FIXED_IO_ps_srstb (FIXED_IO_ps_srstb),
  .FIXED_IO_ddr_vrn  (FIXED_IO_ddr_vrn ),
  .FIXED_IO_ddr_vrp  (FIXED_IO_ddr_vrp ),
  // DDR
  .DDR_addr          (DDR_addr         ),
  .DDR_ba            (DDR_ba           ),
  .DDR_cas_n         (DDR_cas_n        ),
  .DDR_ck_n          (DDR_ck_n         ),
  .DDR_ck_p          (DDR_ck_p         ),
  .DDR_cke           (DDR_cke          ),
  .DDR_cs_n          (DDR_cs_n         ),
  .DDR_dm            (DDR_dm           ),
  .DDR_dq            (DDR_dq           ),
  .DDR_dqs_n         (DDR_dqs_n        ),
  .DDR_dqs_p         (DDR_dqs_p        ),
  .DDR_odt           (DDR_odt          ),
  .DDR_ras_n         (DDR_ras_n        ),
  .DDR_reset_n       (DDR_reset_n      ),
  .DDR_we_n          (DDR_we_n         ),
  // FCLKs
  .FCLK_CLK0         (fclk_clk[0]      ),
  .FCLK_CLK1         (fclk_clk[1]      ),
  .FCLK_CLK2         (fclk_clk[2]      ),
  .FCLK_CLK3         (fclk_clk[3]      ),
  .FCLK_RESET0_N     (fclk_rstn[0]     ),
  .FCLK_RESET1_N     (fclk_rstn[1]     ),
  .FCLK_RESET2_N     (fclk_rstn[2]     ),
  .FCLK_RESET3_N     (fclk_rstn[3]     ),
//  // XADC
//  .Vaux0_v_n (vinn_i[1]),  .Vaux0_v_p (vinp_i[1]),
//  .Vaux1_v_n (vinn_i[2]),  .Vaux1_v_p (vinp_i[2]),
//  .Vaux8_v_n (vinn_i[0]),  .Vaux8_v_p (vinp_i[0]),
//  .Vaux9_v_n (vinn_i[3]),  .Vaux9_v_p (vinp_i[3]),
//  .Vp_Vn_v_n (vinn_i[4]),  .Vp_Vn_v_p (vinp_i[4]),
  // GP0
  .M_AXI_GP0_ACLK    (axi_gp.ACLK   ),
//  .M_AXI_GP0_ARESETn (axi_gp.ARESETn),
  .M_AXI_GP0_arvalid (axi_gp.ARVALID),
  .M_AXI_GP0_awvalid (axi_gp.AWVALID),
  .M_AXI_GP0_bready  (axi_gp.BREADY ),
  .M_AXI_GP0_rready  (axi_gp.RREADY ),
  .M_AXI_GP0_wlast   (axi_gp.WLAST  ),
  .M_AXI_GP0_wvalid  (axi_gp.WVALID ),
  .M_AXI_GP0_arid    (axi_gp.ARID   ),
  .M_AXI_GP0_awid    (axi_gp.AWID   ),
  .M_AXI_GP0_wid     (axi_gp.WID    ),
  .M_AXI_GP0_arburst (axi_gp.ARBURST),
  .M_AXI_GP0_arlock  (axi_gp.ARLOCK ),
  .M_AXI_GP0_arsize  (axi_gp.ARSIZE ),
  .M_AXI_GP0_awburst (axi_gp.AWBURST),
  .M_AXI_GP0_awlock  (axi_gp.AWLOCK ),
  .M_AXI_GP0_awsize  (axi_gp.AWSIZE ),
  .M_AXI_GP0_arprot  (axi_gp.ARPROT ),
  .M_AXI_GP0_awprot  (axi_gp.AWPROT ),
  .M_AXI_GP0_araddr  (axi_gp.ARADDR ),
  .M_AXI_GP0_awaddr  (axi_gp.AWADDR ),
  .M_AXI_GP0_wdata   (axi_gp.WDATA  ),
  .M_AXI_GP0_arcache (axi_gp.ARCACHE),
  .M_AXI_GP0_arlen   (axi_gp.ARLEN  ),
  .M_AXI_GP0_arqos   (axi_gp.ARQOS  ),
  .M_AXI_GP0_awcache (axi_gp.AWCACHE),
  .M_AXI_GP0_awlen   (axi_gp.AWLEN  ),
  .M_AXI_GP0_awqos   (axi_gp.AWQOS  ),
  .M_AXI_GP0_wstrb   (axi_gp.WSTRB  ),
  .M_AXI_GP0_arready (axi_gp.ARREADY),
  .M_AXI_GP0_awready (axi_gp.AWREADY),
  .M_AXI_GP0_bvalid  (axi_gp.BVALID ),
  .M_AXI_GP0_rlast   (axi_gp.RLAST  ),
  .M_AXI_GP0_rvalid  (axi_gp.RVALID ),
  .M_AXI_GP0_wready  (axi_gp.WREADY ),
  .M_AXI_GP0_bid     (axi_gp.BID    ),
  .M_AXI_GP0_rid     (axi_gp.RID    ),
  .M_AXI_GP0_bresp   (axi_gp.BRESP  ),
  .M_AXI_GP0_rresp   (axi_gp.RRESP  ),
  .M_AXI_GP0_rdata   (axi_gp.RDATA  ),
  // AXI4-Lite
  .M_AXI4_LITE_0_araddr  (axi4_lite.ARADDR ),
  .M_AXI4_LITE_0_arprot  (axi4_lite.ARPROT ),
  .M_AXI4_LITE_0_arready (axi4_lite.ARREADY),
  .M_AXI4_LITE_0_arvalid (axi4_lite.ARVALID),
  .M_AXI4_LITE_0_awaddr  (axi4_lite.AWADDR ),
  .M_AXI4_LITE_0_awprot  (axi4_lite.AWPROT ),
  .M_AXI4_LITE_0_awready (axi4_lite.AWREADY),
  .M_AXI4_LITE_0_awvalid (axi4_lite.AWVALID),
  .M_AXI4_LITE_0_bready  (axi4_lite.BREADY ),
  .M_AXI4_LITE_0_bresp   (axi4_lite.BRESP  ),
  .M_AXI4_LITE_0_bvalid  (axi4_lite.BVALID ),
  .M_AXI4_LITE_0_rdata   (axi4_lite.RDATA  ),
  .M_AXI4_LITE_0_rready  (axi4_lite.RREADY ),
  .M_AXI4_LITE_0_rresp   (axi4_lite.RRESP  ),
  .M_AXI4_LITE_0_rvalid  (axi4_lite.RVALID ),
  .M_AXI4_LITE_0_wdata   (axi4_lite.WDATA  ),
  .M_AXI4_LITE_0_wready  (axi4_lite.WREADY ),
  .M_AXI4_LITE_0_wstrb   (axi4_lite.WSTRB  ),
  .M_AXI4_LITE_0_wvalid  (axi4_lite.WVALID )
  // AXI-4 streaming interfaces
//  .S_AXI_STR1_aclk   (sti[1].clk ),  .S_AXI_STR0_aclk   (sti[0].clk ),
//  .S_AXI_STR1_arstn  (sti[1].rstn),  .S_AXI_STR0_arstn  (sti[0].rstn),
//  .S_AXI_STR1_tdata  (sti[1].dat ),  .S_AXI_STR0_tdata  (sti[0].dat ),
//  .S_AXI_STR1_tkeep  ('1         ),  .S_AXI_STR0_tkeep  ('1         ),
//  .S_AXI_STR1_tlast  (sti[1].lst ),  .S_AXI_STR0_tlast  (sti[0].lst ),
//  .S_AXI_STR1_tready (sti[1].rdy ),  .S_AXI_STR0_tready (sti[0].rdy ),
//  .S_AXI_STR1_tvalid (sti[1].vld ),  .S_AXI_STR0_tvalid (sti[0].vld )
);

assign sti[0].rdy = 1'b1;
assign sti[1].rdy = 1'b1;

// since the PS GP0 port is AXI3 and the local bus is AXI4
assign axi_gp.AWREGION = '0;
assign axi_gp.ARREGION = '0;

endmodule
